`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/12/05 21:37:02
// Design Name: 
// Module Name: RF
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module RF(input clk,//��Ƶ�����ʱ�ӣ�ʵ������ʱ��Ū��CPU_clk
input rst,
input RFWr,//mem2reg��дʹ���ź�
input [15:0]sw_i,
input [4:0]A1,A2,A3,//�ڼ����Ĵ���,sw_i��11��8ָ���Ĵ�����
input [31:0]WD,//write data��sw_i��7��4����д������
output [31:0]RD1,RD2
    );
reg [31:0] rf[31:0];//����32���Ĵ���
always@(posedge clk or negedge rst)
begin
    if(!rst)
    begin
    for(integer i=0;i<8;i=i+1)
    begin
    rf[i]=i;
    end
    end
    else begin
    if(RFWr&&(!sw_i[1]))//�ǵ���ģʽ������д���ź���Ч���Ĵ���ֵ���Ա��޸�
    begin 
        rf[A3]=WD;//�Ĵ���A3��ֵ��Ϊ�������ֵ,���з�����
    end
    end
end
//integer i;
//always@(posedge clk or negedge rst)begin
//if(!rst)
//begin
//for(i=0;i<6;i=i+1)
//begin rf[i]=i;end
//end
//else begin
//if(RFWr&&(!sw_i[1]))//�ǵ���ģʽ������д���ź���Ч���Ĵ���ֵ���Ա��޸�
//begin 
//    rf[A3]=WD;//�Ĵ���A3��ֵ��Ϊ�������ֵ,���з�����
//end
//end
//end
assign RD1=(A1!=0)?rf[A1]:0;
assign RD2=(A2!=0)?rf[A2]:0;//������Ĵ�������0�żĴ����������ԭ����ֵ
endmodule
