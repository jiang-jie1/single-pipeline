`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/12/07 20:10:30
// Design Name: 
// Module Name: ALU
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

//A��BΪ����������������ALUopѡ�����ʲô���㣬CΪ�������Ľ����ZeroΪ�����Ƿ����
module ALU(input signed[31:0] A,B,input[4:0] ALUOp,output reg signed[31:0] C,output reg Zero);
//�������
//`define ALUOp_add 5'b00001
//`define ALUOp_sub 5'b00000//��һ��ʵ��
`define ALUOp_add 5'b00001
`define ALUOp_sub 5'b00010//�ڶ���ʵ��

always@(*)
begin
case(ALUOp)
`ALUOp_add:C=A+B;
`ALUOp_sub:C=A-B;
endcase
Zero=(C==0)?1:0;
end
endmodule
