`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/12/07 22:18:32
// Design Name: 
// Module Name: DM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

//DMWrд�źţ�6λ��ַ��32λ���ݣ�DMType�ĵ�����3�֣�sw_i[4:3],��������Ǵ�DM�����ַ�ó�������
module DM(input clk,input DMWr,input[5:0]addr,input [31:0]din,input [2:0]DMType,output reg [31:0]dout   );
reg [7:0]dmem[6:0];//��ά���飬7��8λ��
//��������
`define dm_byte 3'b011
`define dm_halfword 3'b001
`define dm_word 3'b000

//��ʼ��128����Ԫ
initial begin
dmem[0]=8'b00000000;
dmem[1]=8'b00000001;
dmem[2]=8'b00000010;
dmem[3]=8'b00000011;
dmem[4]=8'b00000100;
dmem[5]=8'b00000101;
dmem[6]=8'b00000110;
end
always@(posedge clk)
begin
if(DMWr==1'b1)//д�ź�Ϊ1,���������ַ�������������
begin
case(DMType)
`dm_byte:dmem[addr]<=din[7:0];//��ַ��64�֣�����64���ڴ浥Ԫ��ÿ���ڴ浥Ԫ��8λ
`dm_halfword:begin dmem[addr]<=din[7:0];dmem[addr+1]<=din[15:8]; end
`dm_word:begin dmem[addr]<=din[7:0];dmem[addr+1]<=din[15:8];dmem[addr+2]<=din[23:16];dmem[addr+3]<=din[31:24];end
endcase
end
end

always@(*)
begin
case(DMType)
`dm_byte:dout={{24{dmem[addr][7]}},dmem[addr][7:0]};//24{dmem[addr][7]}��ζ�Ű�dmem[addr][7]����24�Σ�Ҳ���Ƿ�����չ������
`dm_halfword:dout={{16{dmem[addr+1][7]}},dmem[addr+1][7:0],dmem[addr][7:0]};
`dm_word:dout={{16{dmem[addr+1][7]}},dmem[addr+1][7:0],dmem[addr][7:0]};
endcase
end
endmodule
